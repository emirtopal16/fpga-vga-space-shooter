module seven_segment(input [3:0]  N,
                     output [6:0] disp);

   assign disp = (N == 4'h0) ? (7'b1000000) :
                 (N == 4'h1) ? (7'b1111001) :
                 (N == 4'h2) ? (7'b0100100) :
                 (N == 4'h3) ? (7'b0110000) :
                 (N == 4'h4) ? (7'b0011001) :
                 (N == 4'h5) ? (7'b0010010) :
                 (N == 4'h6) ? (7'b0000010) :
                 (N == 4'h7) ? (7'b1111000) :
                 (N == 4'h8) ? (7'b0000000) :
                 (N == 4'h9) ? (7'b0010000) :
                 (N == 4'hA) ? (7'b0001000) :
                 (N == 4'hB) ? (7'b0000011) :
                 (N == 4'hC) ? (7'b1000110) :
                 (N == 4'hD) ? (7'b0100001) :
                 (N == 4'hE) ? (7'b0000110) :
                 (N == 4'hF) ? (7'b0001110) : (7'b1111111);

endmodule // seven_segment
